
// Efinity Top-level template
// Version: 2023.1.150.1.5
// Date: 2023-11-13 18:00

// Copyright (C) 2017 - 2023 Efinix Inc. All rights reserved.

// This file may be used as a starting point for Efinity synthesis top-level target.
// The port list here matches what is expected by Efinity constraint files generated
// by the Efinity Interface Designer.

// To use this:
//     #1)  Save this file with a different name to a different directory, where source files are kept.
//              Example: you may wish to save as F:\FPGA_PRJ\YLS\Nearest_900p_108MHZ_v5_1\efinity_project\DDR3_MC.v
//     #2)  Add the newly saved file into Efinity project as design file
//     #3)  Edit the top level entity in Efinity project to:  DDR3_MC
//     #4)  Insert design content.


module DDR3_MC
(
  input inf_in,
  input nrst,
  input DDR3_PLL_CLKOUT4,
  input DDR3_PLL_LOCK,
  input SYS_PLL_LOCK,
  input hdmi_rx_pll_LOCKED,
  input hdmi_tx_pll_LOCKED,
  input twd_clk,
  input tac_clk,
  input tdqss_clk,
  input sys_clk,
  input clk_10m,
  input core_clk,
  input rxc1,
  input rxc,
  input pll_inst4_CLKOUT0,
  input hdmi_tx_fast_clk,
  input clk_25m,
  input hdmi_rx_fast_clk,
  input i_sysclk_div_2,
  input hdmi_rx_slow_clk,
  input fb,
  input clk_125m,
  input hdmi_tx_4x_clk,
  input osc_clk,
  input hdmi_tx_slow_clk,
  input jtag_inst1_CAPTURE,
  input jtag_inst1_DRCK,
  input jtag_inst1_RESET,
  input jtag_inst1_RUNTEST,
  input jtag_inst1_SEL,
  input jtag_inst1_SHIFT,
  input jtag_inst1_TCK,
  input jtag_inst1_TDI,
  input jtag_inst1_TMS,
  input jtag_inst1_UPDATE,
  input hdmi_rx_clk_RX_DATA,
  input [9:0] hdmi_rx_d0_RX_DATA,
  input [9:0] hdmi_rx_d1_RX_DATA,
  input [9:0] hdmi_rx_d2_RX_DATA,
  input FPGA_HDMI_SCL_IN,
  input FPGA_HDMI_SDA_IN,
  input HDMI_5V_N,
  input [15:0] i_dq_hi,
  input [15:0] i_dq_lo,
  input [1:0] i_dqs_hi,
  input [1:0] i_dqs_lo,
  input hdmi_tx_clk,
  input mdio_i,
  input mdio_io1_IN,
  input rx_dv_HI,
  input rx_dv_LO,
  input rx_dv1_HI,
  input rx_dv1_LO,
  input [3:0] rxd1_HI,
  input [3:0] rxd1_LO,
  input [3:0] rxd_hi_i,
  input [3:0] rxd_lo_i,
  input uart_rx,
  output LCD_POWER,
  output [1:0] b_led,
  output beep,
  output o_lcd_rstn,
  output phy_rst_n,
  output phy_rst_n1,
  output DDR3_PLL_RSTN,
  output [2:0] shift,
  output shift_ena,
  output [4:0] shift_sel,
  output SYS_PLL_RSTN,
  output hdmi_rx_pll_RSTN,
  output hdmi_tx_pll_RSTN,
  output jtag_inst1_TDO,
  output hdmi_rx_clk_RX_ENA,
  output hdmi_rx_d0_RX_RST,
  output hdmi_rx_d0_RX_ENA,
  output hdmi_rx_d1_RX_RST,
  output hdmi_rx_d1_RX_ENA,
  output hdmi_rx_d2_RX_RST,
  output hdmi_rx_d2_RX_ENA,
  output tmds_tx_clk_TX_OE,
  output [9:0] tmds_tx_clk_TX_DATA,
  output tmds_tx_clk_TX_RST,
  output tmds_tx_data0_TX_OE,
  output [9:0] tmds_tx_data0_TX_DATA,
  output tmds_tx_data0_TX_RST,
  output tmds_tx_data1_TX_OE,
  output [9:0] tmds_tx_data1_TX_DATA,
  output tmds_tx_data1_TX_RST,
  output tmds_tx_data2_TX_OE,
  output [9:0] tmds_tx_data2_TX_DATA,
  output tmds_tx_data2_TX_RST,
  output FPGA_HDMI_SCL_OUT,
  output FPGA_HDMI_SCL_OE,
  output FPGA_HDMI_SDA_OUT,
  output FPGA_HDMI_SDA_OE,
  output HPD_N,
  output [15:0] addr,
  output [2:0] ba,
  output cas,
  output cke,
  output cs,
  output [1:0] o_dm_hi,
  output [1:0] o_dm_lo,
  output [15:0] o_dq_hi,
  output [15:0] o_dq_lo,
  output [15:0] o_dq_oe,
  output [1:0] o_dqs_hi,
  output [1:0] o_dqs_lo,
  output [1:0] o_dqs_oe,
  output [1:0] o_dqs_n_oe,
  output mdc_o_HI,
  output mdc_o_LO,
  output mdc_o1_HI,
  output mdc_o1_LO,
  output mdio_o,
  output mdio_oe,
  output mdio_io1_OUT,
  output mdio_io1_OE,
  output odt,
  output ras,
  output reset,
  output tx_en_o_HI,
  output tx_en_o_LO,
  output tx_en_o1_HI,
  output tx_en_o1_LO,
  output txc_hi_o,
  output txc_lo_o,
  output txc1_HI,
  output txc1_LO,
  output [3:0] txd1_HI,
  output [3:0] txd1_LO,
  output [3:0] txd_hi_o,
  output [3:0] txd_lo_o,
  output uart_tx,
  output we,
  output osc_en
);


endmodule

